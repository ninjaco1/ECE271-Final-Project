//Counter and comparator
module 