// shift register

//module shift_register8(input logic clk,input logic [7:0] botton, output logic data); 
//	always_latch
//		if(clk) 
//endmodule
