//Top Level

module FinalProject (input logic clk, ltch, data,
							output logic led, motor,
							output logic [6:0]seg);
							
	
							
	//log						
							
							

endmodule
				