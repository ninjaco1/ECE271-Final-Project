//NES decoder

module NesDecoder (input logic nes_clk, nes_latch,
						input logic [7:0] readButtons,
						output logic );