//Top Level